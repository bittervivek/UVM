//create a interface
//remember to decalare clk, coming from top module
//every signal that comes from top module need to declare as input
Interface our_interface(input );
 //input_1/2
logic input_1
logic input_2

//output
Output output_3

endinterface
